class axi_base_txn extends uvm_sequence_item;
  `uvm_object_utils(axi_base_txn)
  function new(string name="axi_base_txn");
    super.new(name);
  endfunction
endclass
