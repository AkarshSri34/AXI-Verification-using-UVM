`include "interface.sv"
`include "transaction.sv"
`include "slave_transaction.sv"
`include "sequence.sv"
`include "sequencer.sv"
`include "slave_sequencer.sv"
`include "driver.sv"
`include "slave_driver.sv"
//`include "monitor.sv"
`include "agent.sv"
`include "slave_agent.sv"
`include "env.sv"
`include "test.sv"
