class axi_slave_txn extends uvm_sequence_item;
  `uvm_object_utils(axi_slave_txn)
  function new(string name="axi_slave_txn");
    super.new(name);
  endfunction
endclass
